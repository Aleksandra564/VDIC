`timescale 1ns/1ps

package mult_pkg;

	`include "tpgen.svh"
	`include "coverage.svh"
	`include "scoreboard.svh"
	`include "testbench.svh"
	
endpackage : mult_pkg
	